//吃到之後消失
//type 表示顏色 
//後續變數只需要輸入相應的角色
//要寫被吃掉的行為(消失)
module treasure(

);
endmodule