module map(
    input clk, 
    input rst, 
    input en, 
    input [2:0] level,
    input [2:0] map,
    input wire [9:0] vga_h, //640 ?{?b?????X?????pixel
    input wire [9:0] vga_v,  //480 ?{?b?????X?????pixel
    inout PS2_DATA, 
    inout PS2_CLK, 
    output wire [16:0] addr, 
    output reg clear
);

    //player player1(...);
    //player player2(...);
    //terrain t1(...); ...
    //mech m1(...); ...
    wire [16:0] menu_addr;
    assign menu_addr = (level == 0) ? (
        (map == 0) ? (
            ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 40 && (vga_v>>1) <= 65) ? (
                ((vga_h >> 1)-150 + ((vga_v >> 1)-39)*320)
            ) : (
                ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 80 && (vga_v>>1) <= 105) ? (
                    ((vga_h >> 1)-150 + ((vga_v >> 1)-79)*320)
                ): (
                    ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 120 && (vga_v>>1) <= 145) ? (
                        ((vga_h >> 1)-150 + ((vga_v >> 1)-119)*320)
                    ) : (
                        ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 160 && (vga_v>>1) <= 185) ? (
                            ((vga_h >> 1)-150 + ((vga_v >> 1)-159)*320)
                        ) : (
                            ((vga_h>>1) >= 148 && (vga_h>>1) <= 170 && (vga_v>>1) >= 200 && (vga_v>>1) <= 225) ? (
                                ((vga_h >> 1)-127 + ((vga_v >> 1)-199)*320)
                            ) : (
                                0
                            )
                        )
                    )
                )
            )
        ) : (
            (map == 1) ? (
                ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 40 && (vga_v>>1) <= 65) ? (
                    ((vga_h >> 1)-150 + ((vga_v >> 1)-39)*320)
                ) : (
                    ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 80 && (vga_v>>1) <= 105) ? (
                        ((vga_h >> 1)-150 + ((vga_v >> 1)-79)*320)
                    ) : (
                        ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 120 && (vga_v>>1) <= 145) ? (
                            ((vga_h >> 1)-150 + ((vga_v >> 1)-119)*320)
                        ) : (
                            ((vga_h>>1) >= 148 && (vga_h>>1) <= 170 && (vga_v>>1) >= 160 && (vga_v>>1) <= 185) ? (
                                ((vga_h >> 1)-127 + ((vga_v >> 1)-159)*320)
                            ) : (
                                ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 200 && (vga_v>>1) <= 225) ? (
                                    ((vga_h >> 1)-150 + ((vga_v >> 1)-199)*320)
                                ) : (
                                    0
                                )
                            )
                        )
                    )
                )
            ) : (
                (map == 2) ? (
                    ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 40 && (vga_v>>1) <= 65) ? (
                        ((vga_h >> 1)-150 + ((vga_v >> 1)-39)*320)
                    ) : (
                        ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 80 && (vga_v>>1) <= 105) ? (
                            ((vga_h >> 1)-150 + ((vga_v >> 1)-79)*320)
                        ) : (
                            ((vga_h>>1) >= 148 && (vga_h>>1) <= 170 && (vga_v>>1) >= 120 && (vga_v>>1) <= 145) ? (
                                ((vga_h >> 1)-127 + ((vga_v >> 1)-119)*320)
                            ) : (
                                ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 160 && (vga_v>>1) <= 185) ? (
                                    ((vga_h >> 1)-150 + ((vga_v >> 1)-159)*320)
                                ) : (
                                    ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 200 && (vga_v>>1) <= 225) ? (
                                        ((vga_h >> 1)-150 + ((vga_v >> 1)-199)*320)
                                    ) : (
                                        0
                                    )
                                )
                            )
                        )
                    )
                ) : (
                    (map == 3) ? (
                        ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 40 && (vga_v>>1) <= 65) ? (
                            ((vga_h >> 1)-150 + ((vga_v >> 1)-39)*320)
                        ) : (
                            ((vga_h>>1) >= 148 && (vga_h>>1) <= 170 && (vga_v>>1) >= 80 && (vga_v>>1) <= 105) ? (
                                ((vga_h >> 1)-127 + ((vga_v >> 1)-79)*320)
                            ) : (
                                ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 120 && (vga_v>>1) <= 145) ? (
                                    ((vga_h >> 1)-150 + ((vga_v >> 1)-119)*320)
                                ) : (
                                    ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 160 && (vga_v>>1) <= 185) ? (
                                        ((vga_h >> 1)-150 + ((vga_v >> 1)-159)*320)
                                    ) : (
                                        ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 200 && (vga_v>>1) <= 225) ? (
                                            ((vga_h >> 1)-150 + ((vga_v >> 1)-199)*320)
                                        ) : (
                                            0
                                        )
                                    )
                                )
                            )
                        )
                    ) : (
                        (map == 4) ? (
                            ((vga_h>>1) >= 148 && (vga_h>>1) <= 170 && (vga_v>>1) >= 40 && (vga_v>>1) <= 65) ? (
                                ((vga_h >> 1)-127 + ((vga_v >> 1)-39)*320)
                            ) : (
                                ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 80 && (vga_v>>1) <= 105) ? (
                                    ((vga_h >> 1)-150 + ((vga_v >> 1)-79)*320)
                                ) : (
                                    ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 120 && (vga_v>>1) <= 145) ? (
                                        ((vga_h >> 1)-150 + ((vga_v >> 1)-119)*320)
                                    ) : (
                                        ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 160 && (vga_v>>1) <= 185) ? (
                                            ((vga_h >> 1)-150 + ((vga_v >> 1)-159)*320)
                                        ) : (
                                            ((vga_h>>1) >= 150 && (vga_h>>1) <= 170 && (vga_v>>1) >= 200 && (vga_v>>1) <= 225) ? (
                                                ((vga_h >> 1)-150 + ((vga_v >> 1)-199)*320)
                                            ) : (
                                                0
                                            )
                                        )
                                    )
                                )
                            )
                        ) : (

                        )
                    )
                )
            )
        )
    ) : (
        0
    );

    assign addr = (level == 0) ? menu_addr : 0;

endmodule